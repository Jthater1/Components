* NGSPICE file created from 4-1MUX.ext - technology: sky130B

.subckt x4-1MUX S1 B OUT A D C VSS VDD S2
X0 VSS.t2 S2.t0 x3.x3.Vout VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X1 x3.B.t3 x3.x3.Vout OUT.t2 VSS.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X2 A.t1 S1.t0 x3.A VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X3 C.t1 S1.t1 x3.B.t1 VSS.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X4 C.t0 x2.x3.Vout x3.B.t4 VDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5 A.t0 x1.x3.Vout x3.A VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6 VDD.t2 S2.t1 x3.x3.Vout VDD.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7 x3.A S2.t2 OUT.t1 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X8 B.t0 x1.x3.Vout x3.A VSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X9 VDD.t11 S1.t2 x1.x3.Vout VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X10 x3.A x3.x3.Vout OUT.t3 VDD.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X11 VSS.t5 S1.t3 x2.x3.Vout VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X12 VDD.t9 S1.t4 x2.x3.Vout VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X13 B.t1 S1.t5 x3.A VDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X14 VSS.t11 S1.t6 x1.x3.Vout VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X15 D.t0 x2.x3.Vout x3.B.t5 VSS.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X16 D.t1 S1.t7 x3.B.t2 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X17 x3.B.t0 S2.t3 OUT.t0 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
R0 S2.n0 S2.t1 133.2
R1 S2 S2.t3 133.085
R2 S2.n0 S2.t0 112.76
R3 S2 S2.t2 112.734
R4 S2.n2 S2 13.4173
R5 S2.n4 S2 12.9083
R6 S2.n3 S2 11.2052
R7 S2.n2 S2.n1 9.03988
R8 S2.n3 S2.n2 2.20853
R9 S2.n1 S2.n0 0.80869
R10 S2.n4 S2.n3 0.63912
R11 S2 S2.n4 0.061125
R12 S2.n1 S2 0.056125
R13 VSS.n35 VSS.n34 40832.8
R14 VSS.n64 VSS.n63 32392.6
R15 VSS.n68 VSS.n67 30929.4
R16 VSS.n63 VSS.n36 29592.2
R17 VSS.n69 VSS.n68 21769.5
R18 VSS.n118 VSS.n117 19768.3
R19 VSS.n21 VSS.n20 17682
R20 VSS.n68 VSS.n34 17412.2
R21 VSS.n95 VSS.n45 12334.7
R22 VSS.n22 VSS.n16 11233.1
R23 VSS.n118 VSS.n35 9824.14
R24 VSS.n78 VSS.n50 6854.42
R25 VSS.n20 VSS.n16 5182.22
R26 VSS.n117 VSS.n36 3731.37
R27 VSS.n79 VSS.n78 3033.11
R28 VSS.n105 VSS.n104 2847.63
R29 VSS.n78 VSS.n77 2398.83
R30 VSS.n21 VSS.n5 2333.12
R31 VSS.n79 VSS.n46 2163.27
R32 VSS.t3 VSS.n80 1914.29
R33 VSS.n119 VSS.n33 1582.38
R34 VSS.n116 VSS.n37 1488.48
R35 VSS.n93 VSS.n37 1488.48
R36 VSS.n93 VSS.n38 1488.48
R37 VSS.n116 VSS.n38 1488.48
R38 VSS.n122 VSS.n4 1488.48
R39 VSS.n123 VSS.n4 1488.48
R40 VSS.n123 VSS.n3 1488.48
R41 VSS.n122 VSS.n3 1488.48
R42 VSS.n32 VSS.n6 1488.48
R43 VSS.n32 VSS.n7 1488.48
R44 VSS.n18 VSS.n7 1488.48
R45 VSS.n18 VSS.n6 1488.48
R46 VSS.n70 VSS.n60 1488.48
R47 VSS.n76 VSS.n60 1488.48
R48 VSS.n76 VSS.n61 1488.48
R49 VSS.n70 VSS.n61 1488.48
R50 VSS.n107 VSS.n44 1488.48
R51 VSS.n108 VSS.n44 1488.48
R52 VSS.n108 VSS.n43 1488.48
R53 VSS.n107 VSS.n43 1488.48
R54 VSS.n82 VSS.n58 1488.48
R55 VSS.n84 VSS.n58 1488.48
R56 VSS.n82 VSS.n59 1488.48
R57 VSS.n91 VSS.n51 1488.48
R58 VSS.n91 VSS.n52 1488.48
R59 VSS.n66 VSS.n52 1488.48
R60 VSS.n66 VSS.n51 1488.48
R61 VSS.n24 VSS.n13 1488.48
R62 VSS.n25 VSS.n13 1488.48
R63 VSS.n25 VSS.n12 1488.48
R64 VSS.n24 VSS.n12 1488.48
R65 VSS.n103 VSS.n47 1488.48
R66 VSS.n103 VSS.n48 1488.48
R67 VSS.n97 VSS.n48 1488.48
R68 VSS.n97 VSS.n47 1488.48
R69 VSS.n119 VSS.n118 1460.43
R70 VSS.n22 VSS.n21 1223.71
R71 VSS.n63 VSS.n35 1177.36
R72 VSS.n20 VSS.n15 1091.18
R73 VSS.n67 VSS.n64 1056.86
R74 VSS.t6 VSS.n45 1027.18
R75 VSS.t6 VSS.n105 1027.18
R76 VSS.n119 VSS.n34 968.135
R77 VSS.n69 VSS.t4 859.476
R78 VSS.n77 VSS.t4 859.476
R79 VSS.n83 VSS.n59 841.096
R80 VSS.n95 VSS.n94 804.139
R81 VSS.t7 VSS.n14 788.236
R82 VSS.n80 VSS.n79 600
R83 VSS.n94 VSS.t8 580.888
R84 VSS.t8 VSS.n36 552.71
R85 VSS.n22 VSS.n15 523.529
R86 VSS.n92 VSS.t9 476.637
R87 VSS.n16 VSS.n14 474.045
R88 VSS.t0 VSS.n5 455.642
R89 VSS.t0 VSS.n120 455.642
R90 VSS.n64 VSS.t9 453.517
R91 VSS.n33 VSS.t1 302.05
R92 VSS.n19 VSS.t1 300.836
R93 VSS.t7 VSS.n22 264.707
R94 VSS.n95 VSS.n92 247.212
R95 VSS.n120 VSS.n119 224.421
R96 VSS.t10 VSS.n46 215.017
R97 VSS.n50 VSS.t10 179.417
R98 VSS.n97 VSS.n96 168.362
R99 VSS.n96 VSS.n50 157.06
R100 VSS.n19 VSS.n18 147.269
R101 VSS.n43 VSS.n42 146.25
R102 VSS.n45 VSS.n43 146.25
R103 VSS.n44 VSS.n41 146.25
R104 VSS.n105 VSS.n44 146.25
R105 VSS.n91 VSS.n90 146.25
R106 VSS.n92 VSS.n91 146.25
R107 VSS.n59 VSS.n57 146.25
R108 VSS.n58 VSS.n56 146.25
R109 VSS.n80 VSS.n58 146.25
R110 VSS.n71 VSS.n70 146.25
R111 VSS.n70 VSS.n69 146.25
R112 VSS.n76 VSS.n75 146.25
R113 VSS.n77 VSS.n76 146.25
R114 VSS.n66 VSS.n65 146.25
R115 VSS.n67 VSS.n66 146.25
R116 VSS.n12 VSS.n11 146.25
R117 VSS.n14 VSS.n12 146.25
R118 VSS.n13 VSS.n10 146.25
R119 VSS.n15 VSS.n13 146.25
R120 VSS.n18 VSS.n17 146.25
R121 VSS.n32 VSS.n31 146.25
R122 VSS.n33 VSS.n32 146.25
R123 VSS.n3 VSS.n2 146.25
R124 VSS.n5 VSS.n3 146.25
R125 VSS.n4 VSS.n1 146.25
R126 VSS.n120 VSS.n4 146.25
R127 VSS.n116 VSS.n115 146.25
R128 VSS.n117 VSS.n116 146.25
R129 VSS.n93 VSS.n40 146.25
R130 VSS.n94 VSS.n93 146.25
R131 VSS.n98 VSS.n97 146.25
R132 VSS.n103 VSS.n102 146.25
R133 VSS.n104 VSS.n103 146.25
R134 VSS.n20 VSS.n19 145.845
R135 VSS.n96 VSS.n95 145.835
R136 VSS.n73 VSS.t5 119.695
R137 VSS.n29 VSS.t2 119.695
R138 VSS.n100 VSS.t11 119.695
R139 VSS.n107 VSS.n106 97.5005
R140 VSS.t6 VSS.n107 97.5005
R141 VSS.n109 VSS.n108 97.5005
R142 VSS.n108 VSS.t6 97.5005
R143 VSS.n53 VSS.n51 97.5005
R144 VSS.n51 VSS.t9 97.5005
R145 VSS.n54 VSS.n52 97.5005
R146 VSS.n52 VSS.t9 97.5005
R147 VSS.n82 VSS.n81 97.5005
R148 VSS.t3 VSS.n82 97.5005
R149 VSS.n85 VSS.n84 97.5005
R150 VSS.n72 VSS.n61 97.5005
R151 VSS.n61 VSS.t4 97.5005
R152 VSS.n62 VSS.n60 97.5005
R153 VSS.n60 VSS.t4 97.5005
R154 VSS.n24 VSS.n23 97.5005
R155 VSS.t7 VSS.n24 97.5005
R156 VSS.n26 VSS.n25 97.5005
R157 VSS.n25 VSS.t7 97.5005
R158 VSS.n8 VSS.n6 97.5005
R159 VSS.n6 VSS.t1 97.5005
R160 VSS.n9 VSS.n7 97.5005
R161 VSS.n7 VSS.t1 97.5005
R162 VSS.n122 VSS.n121 97.5005
R163 VSS.t0 VSS.n122 97.5005
R164 VSS.n124 VSS.n123 97.5005
R165 VSS.n123 VSS.t0 97.5005
R166 VSS.n39 VSS.n37 97.5005
R167 VSS.t8 VSS.n37 97.5005
R168 VSS.n114 VSS.n38 97.5005
R169 VSS.t8 VSS.n38 97.5005
R170 VSS.n49 VSS.n47 97.5005
R171 VSS.t10 VSS.n47 97.5005
R172 VSS.n99 VSS.n48 97.5005
R173 VSS.t10 VSS.n48 97.5005
R174 VSS.n72 VSS.n71 95.7785
R175 VSS.n17 VSS.n9 95.7785
R176 VSS.n99 VSS.n98 95.7785
R177 VSS.n115 VSS.n39 94.964
R178 VSS.n106 VSS.n42 94.964
R179 VSS.n65 VSS.n53 94.964
R180 VSS.n81 VSS.n57 94.964
R181 VSS.n121 VSS.n2 94.964
R182 VSS.n23 VSS.n11 94.964
R183 VSS.n71 VSS.n62 94.2726
R184 VSS.n17 VSS.n8 94.2726
R185 VSS.n98 VSS.n49 94.2726
R186 VSS.n115 VSS.n114 89.739
R187 VSS.n109 VSS.n42 89.739
R188 VSS.n65 VSS.n54 89.739
R189 VSS.n85 VSS.n57 89.739
R190 VSS.n124 VSS.n2 89.739
R191 VSS.n26 VSS.n11 89.739
R192 VSS.n104 VSS.n46 82.1945
R193 VSS.n83 VSS.t3 55.0953
R194 VSS.n84 VSS.n83 39.7998
R195 VSS.n75 VSS.n62 32.431
R196 VSS.n31 VSS.n8 32.431
R197 VSS.n102 VSS.n49 32.431
R198 VSS.n40 VSS.n39 31.811
R199 VSS.n106 VSS.n41 31.811
R200 VSS.n90 VSS.n53 31.811
R201 VSS.n81 VSS.n56 31.811
R202 VSS.n121 VSS.n1 31.811
R203 VSS.n23 VSS.n10 31.811
R204 VSS.n74 VSS.n72 27.6091
R205 VSS.n30 VSS.n9 27.6091
R206 VSS.n101 VSS.n99 27.6091
R207 VSS.n114 VSS.n113 25.7297
R208 VSS.n110 VSS.n109 25.7297
R209 VSS.n89 VSS.n54 25.7297
R210 VSS.n86 VSS.n85 25.7297
R211 VSS.n125 VSS.n124 25.7297
R212 VSS.n27 VSS.n26 25.7297
R213 VSS VSS.n112 21.3298
R214 VSS VSS.n88 21.3298
R215 VSS.n28 VSS 21.3298
R216 VSS.n88 VSS 14.5351
R217 VSS VSS.n28 14.5351
R218 VSS.n112 VSS 14.5351
R219 VSS.n75 VSS.n74 4.99776
R220 VSS.n31 VSS.n30 4.99776
R221 VSS.n102 VSS.n101 4.99776
R222 VSS.n113 VSS.n40 4.54104
R223 VSS.n110 VSS.n41 4.54104
R224 VSS.n90 VSS.n89 4.54104
R225 VSS.n86 VSS.n56 4.54104
R226 VSS.n125 VSS.n1 4.54104
R227 VSS.n27 VSS.n10 4.54104
R228 VSS.n55 VSS 2.27041
R229 VSS.n113 VSS 0.884986
R230 VSS.n89 VSS 0.884986
R231 VSS VSS.n27 0.884986
R232 VSS.n74 VSS.n73 0.869897
R233 VSS.n30 VSS.n29 0.869897
R234 VSS.n101 VSS.n100 0.869897
R235 VSS.n87 VSS.n86 0.7755
R236 VSS.n126 VSS.n125 0.7755
R237 VSS.n111 VSS.n110 0.7755
R238 VSS.n88 VSS 0.406092
R239 VSS.n28 VSS 0.406092
R240 VSS.n112 VSS 0.406092
R241 VSS VSS.n126 0.300374
R242 VSS.n87 VSS.n55 0.238499
R243 VSS.n111 VSS.n0 0.236649
R244 VSS VSS.n0 0.1255
R245 VSS VSS.n87 0.109986
R246 VSS.n126 VSS 0.109986
R247 VSS VSS.n111 0.109986
R248 VSS.n55 VSS 0.062375
R249 VSS VSS.n0 0.0617745
R250 VSS.n73 VSS 0.0147241
R251 VSS.n29 VSS 0.0147241
R252 VSS.n100 VSS 0.0147241
R253 OUT.n2 OUT.t0 168.333
R254 OUT.n0 OUT.t3 168.333
R255 OUT.n2 OUT.t2 120.234
R256 OUT.n0 OUT.t1 120.234
R257 OUT.n3 OUT 12.912
R258 OUT OUT.n1 3.20883
R259 OUT.n3 OUT.n2 0.711438
R260 OUT.n1 OUT.n0 0.711438
R261 OUT.n1 OUT 0.063
R262 OUT OUT.n3 0.063
R263 x3.B x3.B.t0 168.339
R264 x3.B x3.B.t2 168.333
R265 x3.B x3.B.t4 168.333
R266 x3.B x3.B.t5 120.234
R267 x3.B x3.B.t1 120.234
R268 x3.B x3.B.t3 120.228
R269 S1.n4 S1.t2 133.2
R270 S1.n0 S1.t4 133.2
R271 S1 S1.t5 133.085
R272 S1 S1.t7 133.085
R273 S1.n4 S1.t6 112.76
R274 S1.n0 S1.t3 112.76
R275 S1 S1.t0 112.734
R276 S1 S1.t1 112.734
R277 S1.n6 S1 13.4173
R278 S1.n2 S1 13.4173
R279 S1.n7 S1 11.2052
R280 S1.n3 S1 11.2052
R281 S1.n6 S1.n5 9.03988
R282 S1.n2 S1.n1 9.03988
R283 S1.n7 S1.n6 2.20853
R284 S1.n3 S1.n2 2.20853
R285 S1.n5 S1.n4 0.80869
R286 S1.n1 S1.n0 0.80869
R287 S1 S1.n7 0.699745
R288 S1 S1.n3 0.699745
R289 S1.n5 S1 0.056125
R290 S1.n1 S1 0.056125
R291 A.n0 A.t0 168.339
R292 A.n0 A.t1 120.228
R293 A.n1 A 10.9131
R294 A.n1 A 3.1255
R295 A A.n0 0.701021
R296 A.n2 A 0.123
R297 A A.n2 0.063
R298 A.n2 A.n1 0.00177551
R299 C.n0 C.t0 168.339
R300 C.n0 C.t1 120.228
R301 C C.n0 0.701021
R302 VDD.n5 VDD.n3 1053.52
R303 VDD.n8 VDD.n2 1053.52
R304 VDD.n28 VDD.n26 1053.52
R305 VDD.n31 VDD.n25 1053.52
R306 VDD.n17 VDD.n15 1053.52
R307 VDD.n20 VDD.n14 1053.52
R308 VDD.n42 VDD.n40 1053.52
R309 VDD.n45 VDD.n39 1053.52
R310 VDD.n65 VDD.n63 1053.52
R311 VDD.n68 VDD.n62 1053.52
R312 VDD.n54 VDD.n52 1053.52
R313 VDD.n57 VDD.n51 1053.52
R314 VDD.n104 VDD.n102 1053.52
R315 VDD.n107 VDD.n101 1053.52
R316 VDD.n91 VDD.n89 1053.52
R317 VDD.n94 VDD.n88 1053.52
R318 VDD.n80 VDD.n78 1053.52
R319 VDD.n83 VDD.n77 1053.52
R320 VDD.n6 VDD.n2 372.587
R321 VDD.n7 VDD.n3 372.587
R322 VDD.n29 VDD.n25 372.587
R323 VDD.n30 VDD.n26 372.587
R324 VDD.n18 VDD.n14 372.587
R325 VDD.n19 VDD.n15 372.587
R326 VDD.n43 VDD.n39 372.587
R327 VDD.n44 VDD.n40 372.587
R328 VDD.n66 VDD.n62 372.587
R329 VDD.n67 VDD.n63 372.587
R330 VDD.n55 VDD.n51 372.587
R331 VDD.n56 VDD.n52 372.587
R332 VDD.n105 VDD.n101 372.587
R333 VDD.n106 VDD.n102 372.587
R334 VDD.n92 VDD.n88 372.587
R335 VDD.n93 VDD.n89 372.587
R336 VDD.n81 VDD.n77 372.587
R337 VDD.n82 VDD.n78 372.587
R338 VDD.n11 VDD.t11 167.714
R339 VDD.n48 VDD.t2 167.714
R340 VDD.n110 VDD.t9 167.714
R341 VDD.n9 VDD.n1 102.305
R342 VDD.n46 VDD.n38 102.305
R343 VDD.n108 VDD.n100 102.305
R344 VDD.n32 VDD.n24 101.602
R345 VDD.n27 VDD.n24 101.602
R346 VDD.n21 VDD.n13 101.602
R347 VDD.n16 VDD.n13 101.602
R348 VDD.n69 VDD.n61 101.602
R349 VDD.n64 VDD.n61 101.602
R350 VDD.n58 VDD.n50 101.602
R351 VDD.n53 VDD.n50 101.602
R352 VDD.n95 VDD.n87 101.602
R353 VDD.n90 VDD.n87 101.602
R354 VDD.n84 VDD.n76 101.602
R355 VDD.n79 VDD.n76 101.602
R356 VDD.n4 VDD.n1 101.165
R357 VDD.n41 VDD.n38 101.165
R358 VDD.n103 VDD.n100 101.165
R359 VDD.n2 VDD.n1 46.2505
R360 VDD.n3 VDD.n0 46.2505
R361 VDD.n25 VDD.n24 46.2505
R362 VDD.n26 VDD.n23 46.2505
R363 VDD.n14 VDD.n13 46.2505
R364 VDD.n15 VDD.n12 46.2505
R365 VDD.n39 VDD.n38 46.2505
R366 VDD.n40 VDD.n37 46.2505
R367 VDD.n62 VDD.n61 46.2505
R368 VDD.n63 VDD.n60 46.2505
R369 VDD.n51 VDD.n50 46.2505
R370 VDD.n52 VDD.n49 46.2505
R371 VDD.n101 VDD.n100 46.2505
R372 VDD.n102 VDD.n99 46.2505
R373 VDD.n88 VDD.n87 46.2505
R374 VDD.n89 VDD.n86 46.2505
R375 VDD.n77 VDD.n76 46.2505
R376 VDD.n78 VDD.n75 46.2505
R377 VDD.n27 VDD.n23 37.2794
R378 VDD.n16 VDD.n12 37.2794
R379 VDD.n64 VDD.n60 37.2794
R380 VDD.n53 VDD.n49 37.2794
R381 VDD.n90 VDD.n86 37.2794
R382 VDD.n79 VDD.n75 37.2794
R383 VDD.n4 VDD.n0 37.2504
R384 VDD.n41 VDD.n37 37.2504
R385 VDD.n103 VDD.n99 37.2504
R386 VDD.n33 VDD.n32 33.2599
R387 VDD.n22 VDD.n21 33.2599
R388 VDD.n70 VDD.n69 33.2599
R389 VDD.n59 VDD.n58 33.2599
R390 VDD.n96 VDD.n95 33.2599
R391 VDD.n85 VDD.n84 33.2599
R392 VDD.n10 VDD.n9 32.9612
R393 VDD.n47 VDD.n46 32.9612
R394 VDD.n109 VDD.n108 32.9612
R395 VDD.n9 VDD.n8 23.1255
R396 VDD.n5 VDD.n4 23.1255
R397 VDD.n32 VDD.n31 23.1255
R398 VDD.n28 VDD.n27 23.1255
R399 VDD.n21 VDD.n20 23.1255
R400 VDD.n17 VDD.n16 23.1255
R401 VDD.n46 VDD.n45 23.1255
R402 VDD.n42 VDD.n41 23.1255
R403 VDD.n69 VDD.n68 23.1255
R404 VDD.n65 VDD.n64 23.1255
R405 VDD.n58 VDD.n57 23.1255
R406 VDD.n54 VDD.n53 23.1255
R407 VDD.n108 VDD.n107 23.1255
R408 VDD.n104 VDD.n103 23.1255
R409 VDD.n95 VDD.n94 23.1255
R410 VDD.n91 VDD.n90 23.1255
R411 VDD.n84 VDD.n83 23.1255
R412 VDD.n80 VDD.n79 23.1255
R413 VDD.n34 VDD 22.9581
R414 VDD.n71 VDD 22.9581
R415 VDD.n97 VDD 22.9581
R416 VDD.n6 VDD.n5 14.6266
R417 VDD.n8 VDD.n7 14.6266
R418 VDD.n29 VDD.n28 14.6266
R419 VDD.n31 VDD.n30 14.6266
R420 VDD.n18 VDD.n17 14.6266
R421 VDD.n20 VDD.n19 14.6266
R422 VDD.n43 VDD.n42 14.6266
R423 VDD.n45 VDD.n44 14.6266
R424 VDD.n66 VDD.n65 14.6266
R425 VDD.n68 VDD.n67 14.6266
R426 VDD.n55 VDD.n54 14.6266
R427 VDD.n57 VDD.n56 14.6266
R428 VDD.n105 VDD.n104 14.6266
R429 VDD.n107 VDD.n106 14.6266
R430 VDD.n92 VDD.n91 14.6266
R431 VDD.n94 VDD.n93 14.6266
R432 VDD.n81 VDD.n80 14.6266
R433 VDD.n83 VDD.n82 14.6266
R434 VDD.n35 VDD.n34 13.9985
R435 VDD.n72 VDD.n71 13.9985
R436 VDD.n98 VDD.n97 13.9985
R437 VDD.n7 VDD.t10 8.17936
R438 VDD.t10 VDD.n6 8.17936
R439 VDD.n30 VDD.t4 8.17936
R440 VDD.t4 VDD.n29 8.17936
R441 VDD.n19 VDD.t7 8.17936
R442 VDD.t7 VDD.n18 8.17936
R443 VDD.n44 VDD.t1 8.17936
R444 VDD.t1 VDD.n43 8.17936
R445 VDD.n67 VDD.t3 8.17936
R446 VDD.t3 VDD.n66 8.17936
R447 VDD.n56 VDD.t0 8.17936
R448 VDD.t0 VDD.n55 8.17936
R449 VDD.n106 VDD.t8 8.17936
R450 VDD.t8 VDD.n105 8.17936
R451 VDD.n93 VDD.t5 8.17936
R452 VDD.t5 VDD.n92 8.17936
R453 VDD.n82 VDD.t6 8.17936
R454 VDD.t6 VDD.n81 8.17936
R455 VDD.n10 VDD.n0 4.12253
R456 VDD.n47 VDD.n37 4.12253
R457 VDD.n109 VDD.n99 4.12253
R458 VDD.n74 VDD.n73 4.10971
R459 VDD.n33 VDD.n23 4.02001
R460 VDD.n22 VDD.n12 4.02001
R461 VDD.n70 VDD.n60 4.02001
R462 VDD.n59 VDD.n49 4.02001
R463 VDD.n96 VDD.n86 4.02001
R464 VDD.n85 VDD.n75 4.02001
R465 VDD VDD.n74 3.95513
R466 VDD.n74 VDD.n36 3.7669
R467 VDD VDD.n33 0.875097
R468 VDD VDD.n22 0.875097
R469 VDD VDD.n70 0.875097
R470 VDD VDD.n59 0.875097
R471 VDD VDD.n96 0.875097
R472 VDD VDD.n85 0.875097
R473 VDD.n11 VDD.n10 0.856491
R474 VDD.n48 VDD.n47 0.856491
R475 VDD.n110 VDD.n109 0.856491
R476 VDD.n34 VDD 0.681406
R477 VDD.n71 VDD 0.681406
R478 VDD.n97 VDD 0.681406
R479 VDD.n98 VDD 0.32041
R480 VDD.n36 VDD.n35 0.31916
R481 VDD.n73 VDD.n72 0.31916
R482 VDD.n36 VDD 0.05675
R483 VDD.n73 VDD 0.05675
R484 VDD.n35 VDD 0.0356331
R485 VDD.n72 VDD 0.0356331
R486 VDD VDD.n98 0.0356331
R487 VDD VDD.n11 0.0119645
R488 VDD VDD.n48 0.0119645
R489 VDD VDD.n110 0.0119645
R490 B.n0 B.t1 168.339
R491 B.n0 B.t0 120.228
R492 B B.n0 0.701021
R493 D.n0 D.t1 168.339
R494 D.n0 D.t0 120.228
R495 D D.n0 0.701021
C0 S1 x1.x3.Vout 0.651f
C1 x3.A x1.x3.Vout 0.378f
C2 A x1.x3.Vout 0.3f
C3 S1 x3.A 0.383f
C4 S1 S2 1.43f
C5 S1 A 0.285f
C6 S2 x3.A 0.288f
C7 A x3.A 0.191f
C8 S1 D 0.399f
C9 S1 x2.x3.Vout 0.655f
C10 D S2 0.00295f
C11 D x2.x3.Vout 0.553f
C12 x3.x3.Vout x3.A 0.3f
C13 x3.x3.Vout S2 0.651f
.ends

