* NGSPICE file created from 2-1MUX.ext - technology: sky130B

.subckt x2-1MUX A OUT B VSS VDD S
X0 A.t1 S.t0 OUT.t3 VSS.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X1 B.t0 x3.Vout OUT.t1 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X2 B.t1 S.t1 OUT.t2 VDD.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3 VSS.t2 S.t2 x3.Vout VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X4 A.t0 x3.Vout OUT.t0 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5 VDD.t2 S.t3 x3.Vout VDD.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
R0 S.n1 S.t3 133.2
R1 S S.t1 133.085
R2 S.n1 S.t2 112.76
R3 S S.t0 112.734
R4 S S.n3 13.4173
R5 S.n0 S 11.2052
R6 S.n3 S.n2 9.03988
R7 S.n3 S.n0 2.20853
R8 S.n2 S.n1 0.80869
R9 S.n0 S 0.699745
R10 S.n2 S 0.056125
R11 OUT.n2 OUT.t2 168.333
R12 OUT.n0 OUT.t0 168.333
R13 OUT.n2 OUT.t1 120.234
R14 OUT.n0 OUT.t3 120.234
R15 OUT.n3 OUT 12.912
R16 OUT OUT.n1 3.20883
R17 OUT.n3 OUT.n2 0.711438
R18 OUT.n1 OUT.n0 0.711438
R19 OUT.n1 OUT 0.063
R20 OUT OUT.n3 0.063
R21 A.n0 A.t0 168.339
R22 A.n0 A.t1 120.228
R23 A A.n0 0.701021
R24 VSS.n20 VSS.n9 17139.7
R25 VSS.n20 VSS.n5 16451.1
R26 VSS.n30 VSS.n29 2522.38
R27 VSS.n32 VSS.n4 1488.48
R28 VSS.n33 VSS.n4 1488.48
R29 VSS.n33 VSS.n3 1488.48
R30 VSS.n32 VSS.n3 1488.48
R31 VSS.n18 VSS.n10 1488.48
R32 VSS.n18 VSS.n11 1488.48
R33 VSS.n13 VSS.n11 1488.48
R34 VSS.n13 VSS.n10 1488.48
R35 VSS.n28 VSS.n6 1488.48
R36 VSS.n28 VSS.n7 1488.48
R37 VSS.n22 VSS.n7 1488.48
R38 VSS.n22 VSS.n6 1488.48
R39 VSS.t3 VSS.n5 1225.78
R40 VSS.n20 VSS.n19 885.25
R41 VSS.t3 VSS.n30 704.366
R42 VSS.n30 VSS.n4 667.664
R43 VSS.t0 VSS.n9 639.48
R44 VSS.n19 VSS.t0 639.48
R45 VSS.n29 VSS.t1 583.763
R46 VSS.n21 VSS.t1 580.894
R47 VSS.n21 VSS.n20 279.166
R48 VSS.n22 VSS.n21 148.656
R49 VSS.n3 VSS.n2 146.25
R50 VSS.n5 VSS.n3 146.25
R51 VSS.n4 VSS.n1 146.25
R52 VSS.n14 VSS.n13 146.25
R53 VSS.n13 VSS.n9 146.25
R54 VSS.n18 VSS.n17 146.25
R55 VSS.n19 VSS.n18 146.25
R56 VSS.n23 VSS.n22 146.25
R57 VSS.n28 VSS.n27 146.25
R58 VSS.n29 VSS.n28 146.25
R59 VSS.n25 VSS.t2 119.695
R60 VSS.n32 VSS.n31 97.5005
R61 VSS.t3 VSS.n32 97.5005
R62 VSS.n34 VSS.n33 97.5005
R63 VSS.n33 VSS.t3 97.5005
R64 VSS.n12 VSS.n10 97.5005
R65 VSS.n10 VSS.t0 97.5005
R66 VSS.n15 VSS.n11 97.5005
R67 VSS.n11 VSS.t0 97.5005
R68 VSS.n8 VSS.n6 97.5005
R69 VSS.n6 VSS.t1 97.5005
R70 VSS.n24 VSS.n7 97.5005
R71 VSS.n7 VSS.t1 97.5005
R72 VSS.n24 VSS.n23 95.7785
R73 VSS.n31 VSS.n2 94.964
R74 VSS.n14 VSS.n12 94.964
R75 VSS.n23 VSS.n8 94.2726
R76 VSS.n34 VSS.n2 89.739
R77 VSS.n15 VSS.n14 89.739
R78 VSS.n27 VSS.n8 32.431
R79 VSS.n31 VSS.n1 31.811
R80 VSS.n17 VSS.n12 31.811
R81 VSS.n26 VSS.n24 27.6091
R82 VSS.n35 VSS.n34 25.7297
R83 VSS.n16 VSS.n15 25.7297
R84 VSS VSS.n0 21.3298
R85 VSS VSS.n0 14.5351
R86 VSS.n27 VSS.n26 4.99776
R87 VSS.n35 VSS.n1 4.54104
R88 VSS.n17 VSS.n16 4.54104
R89 VSS.n16 VSS 0.884986
R90 VSS.n26 VSS.n25 0.869897
R91 VSS.n36 VSS.n35 0.7755
R92 VSS VSS.n0 0.406092
R93 VSS.n36 VSS 0.300374
R94 VSS VSS.n36 0.109986
R95 VSS.n25 VSS 0.0147241
R96 B.n0 B.t1 168.339
R97 B.n0 B.t0 120.228
R98 B B.n0 0.701021
R99 VDD.n29 VDD.n27 1053.52
R100 VDD.n32 VDD.n26 1053.52
R101 VDD.n16 VDD.n14 1053.52
R102 VDD.n19 VDD.n13 1053.52
R103 VDD.n5 VDD.n3 1053.52
R104 VDD.n8 VDD.n2 1053.52
R105 VDD.n30 VDD.n26 372.587
R106 VDD.n31 VDD.n27 372.587
R107 VDD.n17 VDD.n13 372.587
R108 VDD.n18 VDD.n14 372.587
R109 VDD.n6 VDD.n2 372.587
R110 VDD.n7 VDD.n3 372.587
R111 VDD.n35 VDD.t2 167.714
R112 VDD.n33 VDD.n25 102.305
R113 VDD.n20 VDD.n12 101.602
R114 VDD.n15 VDD.n12 101.602
R115 VDD.n9 VDD.n1 101.602
R116 VDD.n4 VDD.n1 101.602
R117 VDD.n28 VDD.n25 101.165
R118 VDD.n26 VDD.n25 46.2505
R119 VDD.n27 VDD.n24 46.2505
R120 VDD.n13 VDD.n12 46.2505
R121 VDD.n14 VDD.n11 46.2505
R122 VDD.n2 VDD.n1 46.2505
R123 VDD.n3 VDD.n0 46.2505
R124 VDD.n15 VDD.n11 37.2794
R125 VDD.n4 VDD.n0 37.2794
R126 VDD.n28 VDD.n24 37.2504
R127 VDD.n21 VDD.n20 33.2599
R128 VDD.n10 VDD.n9 33.2599
R129 VDD.n34 VDD.n33 32.9612
R130 VDD.n33 VDD.n32 23.1255
R131 VDD.n29 VDD.n28 23.1255
R132 VDD.n20 VDD.n19 23.1255
R133 VDD.n16 VDD.n15 23.1255
R134 VDD.n9 VDD.n8 23.1255
R135 VDD.n5 VDD.n4 23.1255
R136 VDD.n22 VDD 22.9581
R137 VDD.n30 VDD.n29 14.6266
R138 VDD.n32 VDD.n31 14.6266
R139 VDD.n17 VDD.n16 14.6266
R140 VDD.n19 VDD.n18 14.6266
R141 VDD.n6 VDD.n5 14.6266
R142 VDD.n8 VDD.n7 14.6266
R143 VDD.n23 VDD.n22 13.9985
R144 VDD.n31 VDD.t1 8.17936
R145 VDD.t1 VDD.n30 8.17936
R146 VDD.n18 VDD.t0 8.17936
R147 VDD.t0 VDD.n17 8.17936
R148 VDD.n7 VDD.t3 8.17936
R149 VDD.t3 VDD.n6 8.17936
R150 VDD.n34 VDD.n24 4.12253
R151 VDD.n21 VDD.n11 4.02001
R152 VDD.n10 VDD.n0 4.02001
R153 VDD VDD.n21 0.875097
R154 VDD VDD.n10 0.875097
R155 VDD.n35 VDD.n34 0.856491
R156 VDD.n22 VDD 0.681406
R157 VDD.n23 VDD 0.37541
R158 VDD VDD.n23 0.0356331
R159 VDD VDD.n35 0.0119645
C0 B VDD 0.646f
C1 B x3.Vout 0.553f
C2 B OUT 0.206f
C3 B A 0.253f
C4 x3.Vout VDD 1.3f
C5 B S 0.392f
C6 OUT VDD 1.14f
C7 A VDD 0.217f
C8 OUT x3.Vout 0.378f
C9 A x3.Vout 0.3f
C10 S VDD 2.12f
C11 OUT A 0.191f
C12 S x3.Vout 0.651f
C13 OUT S 0.367f
C14 A S 0.285f
.ends

