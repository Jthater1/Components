* NGSPICE file created from TransmissionGate.ext - technology: sky130B

.subckt TransmissionGate Out In SP VDD VSS SN
X0 Out.t1 SP.t0 In.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1 Out.t0 SN.t0 In.t0 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
R0 SP SP.t0 133.21
R1 In.n0 In.t1 168.339
R2 In.n0 In.t0 120.228
R3 In In.n0 0.826021
R4 Out.n0 Out.t1 168.333
R5 Out.n0 Out.t0 120.234
R6 Out Out.n0 0.773938
R7 VDD.n8 VDD.n7 1053.52
R8 VDD.n5 VDD.n3 1053.52
R9 VDD.n3 VDD.n2 194.792
R10 VDD.n7 VDD.n6 194.792
R11 VDD.n4 VDD.n1 101.602
R12 VDD.n4 VDD.n0 101.602
R13 VDD.n5 VDD.n4 46.2505
R14 VDD.n9 VDD.n8 46.2505
R15 VDD.n9 VDD.n1 37.2794
R16 VDD.n8 VDD.n2 36.1142
R17 VDD.n6 VDD.n5 36.1142
R18 VDD.n10 VDD.n0 33.2599
R19 VDD.n7 VDD.n1 23.1255
R20 VDD.n3 VDD.n0 23.1255
R21 VDD.n6 VDD.t0 8.55241
R22 VDD.t0 VDD.n2 8.55241
R23 VDD.n10 VDD.n9 4.02001
R24 VDD VDD.n10 0.955742
R25 SN SN.t0 112.859
R26 VSS.n6 VSS.n2 1488.48
R27 VSS.n6 VSS.n3 1488.48
R28 VSS.n7 VSS.n3 1488.48
R29 VSS.n7 VSS.n2 1488.48
R30 VSS.n4 VSS.n2 993.766
R31 VSS.n4 VSS.n3 993.766
R32 VSS.n6 VSS.n5 146.25
R33 VSS.t0 VSS.n6 146.25
R34 VSS.n8 VSS.n7 146.25
R35 VSS.n7 VSS.t0 146.25
R36 VSS.n2 VSS.n0 97.5005
R37 VSS.n3 VSS.n1 97.5005
R38 VSS.n5 VSS.n1 94.964
R39 VSS.n5 VSS.n0 89.739
R40 VSS.n8 VSS.n1 31.811
R41 VSS.n9 VSS.n0 25.7297
R42 VSS.t0 VSS.n4 17.6736
R43 VSS.n9 VSS.n8 4.54104
R44 VSS VSS.n9 0.973638
C0 In Out 0.191f
C1 Out SP 0.215f
C2 Out VDD 0.244f
C3 SN Out 0.128f
C4 In SP 0.281f
C5 In VDD 0.216f
C6 SP VDD 0.602f
C7 SN In 0.213f
C8 SN SP 0.0117f
C9 SN VDD 0.00528f
.ends

