* NGSPICE file created from Inverter.ext - technology: sky130B

.subckt Inverter Vin VDD VSS Vout
X0 Vout.t1 Vin.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X1 Vout.t0 Vin.t1 VDD.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
R0 Vin.n0 Vin.t1 133.161
R1 Vin.n0 Vin.t0 112.722
R2 Vin Vin.n0 0.93369
R3 VSS.n6 VSS.n2 1488.48
R4 VSS.n6 VSS.n3 1488.48
R5 VSS.n7 VSS.n3 1488.48
R6 VSS.n7 VSS.n2 1488.48
R7 VSS.n4 VSS.n2 1047.64
R8 VSS.n4 VSS.n3 1047.64
R9 VSS.n6 VSS.n5 146.25
R10 VSS.t0 VSS.n6 146.25
R11 VSS.n8 VSS.n7 146.25
R12 VSS.n7 VSS.t0 146.25
R13 VSS.n10 VSS.t1 119.695
R14 VSS.n2 VSS.n0 97.5005
R15 VSS.n3 VSS.n1 97.5005
R16 VSS.n5 VSS.n0 95.7785
R17 VSS.n5 VSS.n1 94.2726
R18 VSS.n8 VSS.n1 32.431
R19 VSS.n9 VSS.n0 27.6091
R20 VSS.t0 VSS.n4 20.2778
R21 VSS.n9 VSS.n8 4.99776
R22 VSS.n10 VSS.n9 0.869897
R23 VSS VSS.n10 0.100931
R24 Vout.n0 Vout.t0 168.077
R25 Vout.n0 Vout.t1 119.984
R26 Vout Vout.n0 0.664228
R27 VDD.n8 VDD.n7 1053.52
R28 VDD.n5 VDD.n3 1053.52
R29 VDD.n3 VDD.n2 194.792
R30 VDD.n7 VDD.n6 194.792
R31 VDD.n11 VDD.t1 167.714
R32 VDD.n4 VDD.n0 102.305
R33 VDD.n4 VDD.n1 101.165
R34 VDD.n5 VDD.n4 46.2505
R35 VDD.n9 VDD.n8 46.2505
R36 VDD.n9 VDD.n1 37.2504
R37 VDD.n8 VDD.n2 36.1142
R38 VDD.n6 VDD.n5 36.1142
R39 VDD.n10 VDD.n0 32.9612
R40 VDD.n7 VDD.n1 23.1255
R41 VDD.n3 VDD.n0 23.1255
R42 VDD.n6 VDD.t0 8.55241
R43 VDD.t0 VDD.n2 8.55241
R44 VDD.n10 VDD.n9 4.12253
R45 VDD.n11 VDD.n10 0.856491
R46 VDD VDD.n11 0.085929
C0 Vout Vin 0.537f
C1 VDD Vout 0.3f
C2 VDD Vin 0.652f
.ends

