* NGSPICE file created from Buffer.ext - technology: sky130B

.subckt Buffer VDD VSS Vin Vout
X0 Vout.t0 x1.Vout VDD.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1 x1.Vout Vin.t0 VDD.t3 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2 Vout.t1 x1.Vout VSS.t1 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
X3 x1.Vout Vin.t1 VSS.t3 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.5
R0 VDD.n22 VDD.n4 1053.52
R1 VDD.n19 VDD.n5 1053.52
R2 VDD.n12 VDD.n8 1053.52
R3 VDD.n15 VDD.n14 1053.52
R4 VDD.n20 VDD.n4 194.792
R5 VDD.n21 VDD.n5 194.792
R6 VDD.n15 VDD.n7 194.792
R7 VDD.n13 VDD.n12 194.792
R8 VDD.n1 VDD.t3 167.714
R9 VDD.n0 VDD.t1 167.714
R10 VDD.n18 VDD.n17 103.529
R11 VDD.n11 VDD.n6 102.305
R12 VDD.n17 VDD.n6 101.647
R13 VDD.n18 VDD.n3 101.165
R14 VDD.n9 VDD.n8 46.2505
R15 VDD.n14 VDD.n6 46.2505
R16 VDD.n19 VDD.n18 46.2505
R17 VDD.n23 VDD.n22 46.2505
R18 VDD.n23 VDD.n3 37.2504
R19 VDD.n22 VDD.n21 36.1142
R20 VDD.n20 VDD.n19 36.1142
R21 VDD.n8 VDD.n7 36.1142
R22 VDD.n14 VDD.n13 36.1142
R23 VDD.n11 VDD.n10 32.9612
R24 VDD.n12 VDD.n11 23.1255
R25 VDD.n16 VDD.n15 23.1255
R26 VDD.n16 VDD.n4 23.1255
R27 VDD.n5 VDD.n3 23.1255
R28 VDD.n16 VDD.n2 11.5385
R29 VDD.n13 VDD.t0 8.55241
R30 VDD.t0 VDD.n7 8.55241
R31 VDD.t2 VDD.n20 8.55241
R32 VDD.n21 VDD.t2 8.55241
R33 VDD.n17 VDD.n16 7.5498
R34 VDD.n9 VDD.n2 6.94287
R35 VDD.n10 VDD.n9 4.12253
R36 VDD.n24 VDD.n23 4.12253
R37 VDD.n24 VDD.n2 2.96547
R38 VDD.n10 VDD.n0 0.856491
R39 VDD.n25 VDD.n24 0.7755
R40 VDD VDD.n25 0.18763
R41 VDD VDD.n0 0.085929
R42 VDD.n1 VDD 0.085929
R43 VDD.n25 VDD.n1 0.0814911
R44 Vout.n0 Vout.t0 168.077
R45 Vout.n0 Vout.t1 119.984
R46 Vout Vout.n0 0.664228
R47 Vin.n0 Vin.t0 133.161
R48 Vin.n0 Vin.t1 112.722
R49 Vin Vin.n0 0.93369
R50 VSS.n15 VSS.n5 28929.3
R51 VSS.n15 VSS.n14 28693.5
R52 VSS.n16 VSS.n15 13135.3
R53 VSS.n22 VSS.n2 1488.48
R54 VSS.n22 VSS.n3 1488.48
R55 VSS.n23 VSS.n3 1488.48
R56 VSS.n23 VSS.n2 1488.48
R57 VSS.n13 VSS.n7 1488.48
R58 VSS.n18 VSS.n7 1488.48
R59 VSS.n13 VSS.n8 1488.48
R60 VSS.n18 VSS.n8 1488.48
R61 VSS.n17 VSS.n16 1232.56
R62 VSS.n16 VSS.n4 1232.56
R63 VSS.n14 VSS.t0 990.698
R64 VSS.n17 VSS.t0 990.698
R65 VSS.t2 VSS.n4 990.698
R66 VSS.t2 VSS.n5 990.698
R67 VSS.n7 VSS.n6 146.25
R68 VSS.t0 VSS.n7 146.25
R69 VSS.n9 VSS.n8 146.25
R70 VSS.t0 VSS.n8 146.25
R71 VSS.n22 VSS.n21 146.25
R72 VSS.t2 VSS.n22 146.25
R73 VSS.n24 VSS.n23 146.25
R74 VSS.n23 VSS.t2 146.25
R75 VSS.n10 VSS.t1 119.695
R76 VSS.n27 VSS.t3 119.695
R77 VSS.n13 VSS.n12 97.5005
R78 VSS.n14 VSS.n13 97.5005
R79 VSS.n19 VSS.n18 97.5005
R80 VSS.n18 VSS.n17 97.5005
R81 VSS.n19 VSS.n2 97.5005
R82 VSS.n4 VSS.n2 97.5005
R83 VSS.n3 VSS.n1 97.5005
R84 VSS.n5 VSS.n3 97.5005
R85 VSS.n12 VSS.n6 95.7785
R86 VSS.n21 VSS.n1 94.2726
R87 VSS.n21 VSS.n20 92.2776
R88 VSS.n20 VSS.n6 90.7717
R89 VSS.n24 VSS.n1 32.431
R90 VSS.n12 VSS.n11 27.6091
R91 VSS.n19 VSS.n0 8.94698
R92 VSS.n9 VSS.n0 8.41694
R93 VSS.n20 VSS.n19 5.20613
R94 VSS.n11 VSS.n9 4.99776
R95 VSS.n25 VSS.n24 4.99776
R96 VSS.n25 VSS.n0 3.59502
R97 VSS.n11 VSS.n10 0.869897
R98 VSS.n26 VSS.n25 0.7755
R99 VSS.n26 VSS 0.217741
R100 VSS.n10 VSS 0.100931
R101 VSS VSS.n27 0.100931
R102 VSS.n27 VSS.n26 0.0948966
C0 x1.Vout Vout 0.537f
.ends

